* Parametric Inverter Model using BSIM4
* File: inverter.cir
* Inverter subcircuit
.subckt inverter in out vdd vss tplv=0 tpwv=0 tnlv=0 tnwv=0 tpotv=0 tnotv=0
    * BSIM4 Model Parameters
    .model pmos pmos level=54 version=4.8.2
    + toxe = {2.5e-9 + tpotv}
    + toxp = {2.5e-9 + tpotv}
    + toxm = {2.5e-9 + tpotv}
    + dtox = {0 + tpotv}
    + xl = {0 + tplv}
    + xw = {0 + tpwv}
    * Add other PMOS parameters here if needed

    .model nmos nmos level=54 version=4.8.2
    + toxe = {2.5e-9 + tnotv}
    + toxp = {2.5e-9 + tnotv}
    + toxm = {2.5e-9 + tnotv}
    + dtox = {0 + tnotv}
    + xl = {0 + tnlv}
    + xw = {0 + tnwv}
    * Add other NMOS parameters here if needed

    MP out in vdd vdd pmos w={260n + tpwv} l={130n + tplv}
    MN out in vss vss nmos w={130n + tnwv} l={130n + tnlv}
.ends inverter