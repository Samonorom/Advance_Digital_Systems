.subckt ro_1 enable out vdd vss
X1 enable in feedback vdd vss nand tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X2 feedback n2 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X3 n2 n3 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X4 n3 n4 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X5 n4 n5 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X6 n5 n6 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X7 n6 n7 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X8 n7 n8 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X9 n8 n9 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X10 n9 n10 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X11 n10 n11 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X12 n11 n12 vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
X13 n12 out vdd vss inverter tplv=-4.4587e-09 tpwv=-1.7606e-08 tnlv=1.6976e-09 tnwv=-5.6298e-09 tpotv=-1.0781e-10 tnotv=5.2987e-12
* Feedback connection
* 1 ohm resistor for feedback
Rfeedback out in 1
.ends ro_1
