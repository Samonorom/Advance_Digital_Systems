* Ring Oscillator PUF Simulation

* Include component models
.include inverter.cir
.include nand.cir

* Include ring oscillator subcircuits
.include ring_oscillator_0.cir
.include ring_oscillator_1.cir
.include ring_oscillator_2.cir
.include ring_oscillator_3.cir
.include ring_oscillator_4.cir
.include ring_oscillator_5.cir
.include ring_oscillator_6.cir
.include ring_oscillator_7.cir

* senario variation
* Power supply
Vdd vdd 0 dc 1.2
.temp 13.5

* Enable signal (pulse)
Ven enable 0 PULSE(0 1.2 1n 0.1n 0.1n 98n 100n)

* Instantiate ring oscillators
X0 enable out0 vdd 0 ro_0
X1 enable out1 vdd 0 ro_1
X2 enable out2 vdd 0 ro_2
X3 enable out3 vdd 0 ro_3
X4 enable out4 vdd 0 ro_4
X5 enable out5 vdd 0 ro_5
X6 enable out6 vdd 0 ro_6
X7 enable out7 vdd 0 ro_7

* Simulation control
.control
    * Run transient analysis
    tran 0.1n 10n

    * Plot results
    plot v(enable) v(out0)+vdd  v(out1)+2*vdd v(out2)+3*vdd  v(out3)+4*vdd v(out4)+5*vdd v(out5)+6*vdd v(out6)+7*vdd v(out7)+8*vdd
 

    * Write data to a file
    wrdata ro_puf_simulation.txt v(enable) v(out0) v(out1) v(out2) v(out3) v(out4) v(out5) v(out6) v(out7)
.endc

.end