.subckt ro_4 enable out vdd vss
X1 enable in feedback vdd vss nand tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X2 feedback n2 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X3 n2 n3 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X4 n3 n4 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X5 n4 n5 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X6 n5 n6 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X7 n6 n7 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X8 n7 n8 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X9 n8 n9 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X10 n9 n10 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X11 n10 n11 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X12 n11 n12 vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
X13 n12 out vdd vss inverter tplv=-4.2956e-09 tpwv=8.5774e-09 tnlv=1.0111e-09 tnwv=1.5930e-08 tpotv=-1.8229e-10 tnotv=-1.6309e-11
* Feedback connection
* 1 ohm resistor for feedback
Rfeedback out in 1
.ends ro_4
