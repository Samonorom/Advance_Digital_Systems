.subckt ro_0 enable out vdd vss
X1 enable in feedback vdd vss nand tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X2 feedback n2 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X3 n2 n3 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X4 n3 n4 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X5 n4 n5 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X6 n5 n6 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X7 n6 n7 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X8 n7 n8 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X9 n8 n9 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X10 n9 n10 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X11 n10 n11 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X12 n11 n12 vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
X13 n12 out vdd vss inverter tplv=-4.7599e-09 tpwv=-1.1437e-08 tnlv=1.2984e-08 tnwv=4.7542e-09 tpotv=1.6343e-10 tnotv=5.7088e-11
* Feedback connection
* 1 ohm resistor for feedback
Rfeedback out in 1
.ends ro_0
